`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 17.02.2025 15:09:51
// Design Name: 
// Module Name: full_GF_mult
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module full_GF_mult(
    input [3:0] A,
    input [3:0] B,
    output [3:0] out
    );

reg [3:0] OUT;
assign out = OUT;
//use bit concatenation. 
//e.g. if A = 0011 (3) B = 1010 (10) then {A,B} = 00111010.
//this allows us to select the output based on two different numbers.
//the case looks for 00111010 (AB) and finds the output for that sequence of bits
always@(A, B) begin
    case({A, B})
        8'b00000000: OUT <= 0; // 0 * 0
        8'b00000001: OUT <= 0; // 0 * 1
        8'b00000010: OUT <= 0; // 0 * 2
        8'b00000011: OUT <= 0; // 0 * 3
        8'b00000100: OUT <= 0; // 0 * 4
        8'b00000101: OUT <= 0; // 0 * 5
        8'b00000110: OUT <= 0; // 0 * 6
        8'b00000111: OUT <= 0; // 0 * 7
        8'b00001000: OUT <= 0; // 0 * 8
        8'b00001001: OUT <= 0; // 0 * 9
        8'b00001010: OUT <= 0; // 0 * 10
        8'b00001011: OUT <= 0; // 0 * 11
        8'b00001100: OUT <= 0; // 0 * 12
        8'b00001101: OUT <= 0; // 0 * 13
        8'b00001110: OUT <= 0; // 0 * 14
        8'b00001111: OUT <= 0; // 0 * 15
        8'b00010000: OUT <= 0; // 1 * 0
        8'b00010001: OUT <= 1; // 1 * 1
        8'b00010010: OUT <= 2; // 1 * 2
        8'b00010011: OUT <= 3; // 1 * 3
        8'b00010100: OUT <= 4; // 1 * 4
        8'b00010101: OUT <= 5; // 1 * 5
        8'b00010110: OUT <= 6; // 1 * 6
        8'b00010111: OUT <= 7; // 1 * 7
        8'b00011000: OUT <= 8; // 1 * 8
        8'b00011001: OUT <= 9; // 1 * 9
        8'b00011010: OUT <= 10; // 1 * 10
        8'b00011011: OUT <= 11; // 1 * 11
        8'b00011100: OUT <= 12; // 1 * 12
        8'b00011101: OUT <= 13; // 1 * 13
        8'b00011110: OUT <= 14; // 1 * 14
        8'b00011111: OUT <= 15; // 1 * 15
        8'b00100000: OUT <= 0; // 2 * 0
        8'b00100001: OUT <= 2; // 2 * 1
        8'b00100010: OUT <= 4; // 2 * 2
        8'b00100011: OUT <= 6; // 2 * 3
        8'b00100100: OUT <= 8; // 2 * 4
        8'b00100101: OUT <= 10; // 2 * 5
        8'b00100110: OUT <= 12; // 2 * 6
        8'b00100111: OUT <= 14; // 2 * 7
        8'b00101000: OUT <= 3; // 2 * 8
        8'b00101001: OUT <= 1; // 2 * 9
        8'b00101010: OUT <= 7; // 2 * 10
        8'b00101011: OUT <= 5; // 2 * 11
        8'b00101100: OUT <= 11; // 2 * 12
        8'b00101101: OUT <= 9; // 2 * 13
        8'b00101110: OUT <= 15; // 2 * 14
        8'b00101111: OUT <= 13; // 2 * 15
        8'b00110000: OUT <= 0; // 3 * 0
        8'b00110001: OUT <= 3; // 3 * 1
        8'b00110010: OUT <= 6; // 3 * 2
        8'b00110011: OUT <= 5; // 3 * 3
        8'b00110100: OUT <= 12; // 3 * 4
        8'b00110101: OUT <= 15; // 3 * 5
        8'b00110110: OUT <= 10; // 3 * 6
        8'b00110111: OUT <= 9; // 3 * 7
        8'b00111000: OUT <= 11; // 3 * 8
        8'b00111001: OUT <= 8; // 3 * 9
        8'b00111010: OUT <= 13; // 3 * 10
        8'b00111011: OUT <= 14; // 3 * 11
        8'b00111100: OUT <= 7; // 3 * 12
        8'b00111101: OUT <= 4; // 3 * 13
        8'b00111110: OUT <= 1; // 3 * 14
        8'b00111111: OUT <= 2; // 3 * 15
        8'b01000000: OUT <= 0; // 4 * 0
        8'b01000001: OUT <= 4; // 4 * 1
        8'b01000010: OUT <= 8; // 4 * 2
        8'b01000011: OUT <= 12; // 4 * 3
        8'b01000100: OUT <= 3; // 4 * 4
        8'b01000101: OUT <= 7; // 4 * 5
        8'b01000110: OUT <= 11; // 4 * 6
        8'b01000111: OUT <= 15; // 4 * 7
        8'b01001000: OUT <= 6; // 4 * 8
        8'b01001001: OUT <= 2; // 4 * 9
        8'b01001010: OUT <= 14; // 4 * 10
        8'b01001011: OUT <= 10; // 4 * 11
        8'b01001100: OUT <= 5; // 4 * 12
        8'b01001101: OUT <= 1; // 4 * 13
        8'b01001110: OUT <= 13; // 4 * 14
        8'b01001111: OUT <= 9; // 4 * 15
        8'b01010000: OUT <= 0; // 5 * 0
        8'b01010001: OUT <= 5; // 5 * 1
        8'b01010010: OUT <= 10; // 5 * 2
        8'b01010011: OUT <= 15; // 5 * 3
        8'b01010100: OUT <= 7; // 5 * 4
        8'b01010101: OUT <= 2; // 5 * 5
        8'b01010110: OUT <= 13; // 5 * 6
        8'b01010111: OUT <= 8; // 5 * 7
        8'b01011000: OUT <= 14; // 5 * 8
        8'b01011001: OUT <= 11; // 5 * 9
        8'b01011010: OUT <= 4; // 5 * 10
        8'b01011011: OUT <= 1; // 5 * 11
        8'b01011100: OUT <= 9; // 5 * 12
        8'b01011101: OUT <= 12; // 5 * 13
        8'b01011110: OUT <= 3; // 5 * 14
        8'b01011111: OUT <= 6; // 5 * 15
        8'b01100000: OUT <= 0; // 6 * 0
        8'b01100001: OUT <= 6; // 6 * 1
        8'b01100010: OUT <= 12; // 6 * 2
        8'b01100011: OUT <= 10; // 6 * 3
        8'b01100100: OUT <= 11; // 6 * 4
        8'b01100101: OUT <= 13; // 6 * 5
        8'b01100110: OUT <= 7; // 6 * 6
        8'b01100111: OUT <= 1; // 6 * 7
        8'b01101000: OUT <= 5; // 6 * 8
        8'b01101001: OUT <= 3; // 6 * 9
        8'b01101010: OUT <= 9; // 6 * 10
        8'b01101011: OUT <= 15; // 6 * 11
        8'b01101100: OUT <= 14; // 6 * 12
        8'b01101101: OUT <= 8; // 6 * 13
        8'b01101110: OUT <= 2; // 6 * 14
        8'b01101111: OUT <= 4; // 6 * 15
        8'b01110000: OUT <= 0; // 7 * 0
        8'b01110001: OUT <= 7; // 7 * 1
        8'b01110010: OUT <= 14; // 7 * 2
        8'b01110011: OUT <= 9; // 7 * 3
        8'b01110100: OUT <= 15; // 7 * 4
        8'b01110101: OUT <= 8; // 7 * 5
        8'b01110110: OUT <= 1; // 7 * 6
        8'b01110111: OUT <= 6; // 7 * 7
        8'b01111000: OUT <= 13; // 7 * 8
        8'b01111001: OUT <= 10; // 7 * 9
        8'b01111010: OUT <= 3; // 7 * 10
        8'b01111011: OUT <= 4; // 7 * 11
        8'b01111100: OUT <= 2; // 7 * 12
        8'b01111101: OUT <= 5; // 7 * 13
        8'b01111110: OUT <= 12; // 7 * 14
        8'b01111111: OUT <= 11; // 7 * 15
        8'b10000000: OUT <= 0; // 8 * 0
        8'b10000001: OUT <= 8; // 8 * 1
        8'b10000010: OUT <= 3; // 8 * 2
        8'b10000011: OUT <= 11; // 8 * 3
        8'b10000100: OUT <= 6; // 8 * 4
        8'b10000101: OUT <= 14; // 8 * 5
        8'b10000110: OUT <= 5; // 8 * 6
        8'b10000111: OUT <= 13; // 8 * 7
        8'b10001000: OUT <= 12; // 8 * 8
        8'b10001001: OUT <= 4; // 8 * 9
        8'b10001010: OUT <= 15; // 8 * 10
        8'b10001011: OUT <= 7; // 8 * 11
        8'b10001100: OUT <= 10; // 8 * 12
        8'b10001101: OUT <= 2; // 8 * 13
        8'b10001110: OUT <= 9; // 8 * 14
        8'b10001111: OUT <= 1; // 8 * 15
        8'b10010000: OUT <= 0; // 9 * 0
        8'b10010001: OUT <= 9; // 9 * 1
        8'b10010010: OUT <= 1; // 9 * 2
        8'b10010011: OUT <= 8; // 9 * 3
        8'b10010100: OUT <= 2; // 9 * 4
        8'b10010101: OUT <= 11; // 9 * 5
        8'b10010110: OUT <= 3; // 9 * 6
        8'b10010111: OUT <= 10; // 9 * 7
        8'b10011000: OUT <= 4; // 9 * 8
        8'b10011001: OUT <= 13; // 9 * 9
        8'b10011010: OUT <= 5; // 9 * 10
        8'b10011011: OUT <= 12; // 9 * 11
        8'b10011100: OUT <= 6; // 9 * 12
        8'b10011101: OUT <= 15; // 9 * 13
        8'b10011110: OUT <= 7; // 9 * 14
        8'b10011111: OUT <= 14; // 9 * 15
        8'b10100000: OUT <= 0; // 10 * 0
        8'b10100001: OUT <= 10; // 10 * 1
        8'b10100010: OUT <= 7; // 10 * 2
        8'b10100011: OUT <= 13; // 10 * 3
        8'b10100100: OUT <= 14; // 10 * 4
        8'b10100101: OUT <= 4; // 10 * 5
        8'b10100110: OUT <= 9; // 10 * 6
        8'b10100111: OUT <= 3; // 10 * 7
        8'b10101000: OUT <= 15; // 10 * 8
        8'b10101001: OUT <= 5; // 10 * 9
        8'b10101010: OUT <= 8; // 10 * 10
        8'b10101011: OUT <= 2; // 10 * 11
        8'b10101100: OUT <= 1; // 10 * 12
        8'b10101101: OUT <= 11; // 10 * 13
        8'b10101110: OUT <= 6; // 10 * 14
        8'b10101111: OUT <= 12; // 10 * 15
        8'b10110000: OUT <= 0; // 11 * 0
        8'b10110001: OUT <= 11; // 11 * 1
        8'b10110010: OUT <= 5; // 11 * 2
        8'b10110011: OUT <= 14; // 11 * 3
        8'b10110100: OUT <= 10; // 11 * 4
        8'b10110101: OUT <= 1; // 11 * 5
        8'b10110110: OUT <= 15; // 11 * 6
        8'b10110111: OUT <= 4; // 11 * 7
        8'b10111000: OUT <= 7; // 11 * 8
        8'b10111001: OUT <= 12; // 11 * 9
        8'b10111010: OUT <= 2; // 11 * 10
        8'b10111011: OUT <= 9; // 11 * 11
        8'b10111100: OUT <= 13; // 11 * 12
        8'b10111101: OUT <= 6; // 11 * 13
        8'b10111110: OUT <= 8; // 11 * 14
        8'b10111111: OUT <= 3; // 11 * 15
        8'b11000000: OUT <= 0; // 12 * 0
        8'b11000001: OUT <= 12; // 12 * 1
        8'b11000010: OUT <= 11; // 12 * 2
        8'b11000011: OUT <= 7; // 12 * 3
        8'b11000100: OUT <= 5; // 12 * 4
        8'b11000101: OUT <= 9; // 12 * 5
        8'b11000110: OUT <= 14; // 12 * 6
        8'b11000111: OUT <= 2; // 12 * 7
        8'b11001000: OUT <= 10; // 12 * 8
        8'b11001001: OUT <= 6; // 12 * 9
        8'b11001010: OUT <= 1; // 12 * 10
        8'b11001011: OUT <= 13; // 12 * 11
        8'b11001100: OUT <= 15; // 12 * 12
        8'b11001101: OUT <= 3; // 12 * 13
        8'b11001110: OUT <= 4; // 12 * 14
        8'b11001111: OUT <= 8; // 12 * 15
        8'b11010000: OUT <= 0; // 13 * 0
        8'b11010001: OUT <= 13; // 13 * 1
        8'b11010010: OUT <= 9; // 13 * 2
        8'b11010011: OUT <= 4; // 13 * 3
        8'b11010100: OUT <= 1; // 13 * 4
        8'b11010101: OUT <= 12; // 13 * 5
        8'b11010110: OUT <= 8; // 13 * 6
        8'b11010111: OUT <= 5; // 13 * 7
        8'b11011000: OUT <= 2; // 13 * 8
        8'b11011001: OUT <= 15; // 13 * 9
        8'b11011010: OUT <= 11; // 13 * 10
        8'b11011011: OUT <= 6; // 13 * 11
        8'b11011100: OUT <= 3; // 13 * 12
        8'b11011101: OUT <= 14; // 13 * 13
        8'b11011110: OUT <= 10; // 13 * 14
        8'b11011111: OUT <= 7; // 13 * 15
        8'b11100000: OUT <= 0; // 14 * 0
        8'b11100001: OUT <= 14; // 14 * 1
        8'b11100010: OUT <= 15; // 14 * 2
        8'b11100011: OUT <= 1; // 14 * 3
        8'b11100100: OUT <= 13; // 14 * 4
        8'b11100101: OUT <= 3; // 14 * 5
        8'b11100110: OUT <= 2; // 14 * 6
        8'b11100111: OUT <= 12; // 14 * 7
        8'b11101000: OUT <= 9; // 14 * 8
        8'b11101001: OUT <= 7; // 14 * 9
        8'b11101010: OUT <= 6; // 14 * 10
        8'b11101011: OUT <= 8; // 14 * 11
        8'b11101100: OUT <= 4; // 14 * 12
        8'b11101101: OUT <= 10; // 14 * 13
        8'b11101110: OUT <= 11; // 14 * 14
        8'b11101111: OUT <= 5; // 14 * 15
        8'b11110000: OUT <= 0; // 15 * 0
        8'b11110001: OUT <= 15; // 15 * 1
        8'b11110010: OUT <= 13; // 15 * 2
        8'b11110011: OUT <= 2; // 15 * 3
        8'b11110100: OUT <= 9; // 15 * 4
        8'b11110101: OUT <= 6; // 15 * 5
        8'b11110110: OUT <= 4; // 15 * 6
        8'b11110111: OUT <= 11; // 15 * 7
        8'b11111000: OUT <= 1; // 15 * 8
        8'b11111001: OUT <= 14; // 15 * 9
        8'b11111010: OUT <= 12; // 15 * 10
        8'b11111011: OUT <= 3; // 15 * 11
        8'b11111100: OUT <= 8; // 15 * 12
        8'b11111101: OUT <= 7; // 15 * 13
        8'b11111110: OUT <= 5; // 15 * 14
        8'b11111111: OUT <= 10; // 15 * 15
        default: OUT <= 0;
    endcase
end

endmodule
